
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/11/2021 09:44:35 PM
// Design Name: 
// Module Name: axi_intercon_WR
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module axi_intercon_wr (
    input  wire        clk_i,
    input  wire        rst_ni,
    input  wire  [2:0] i_ifu_arid,
    input  wire [31:0] i_ifu_araddr,
    input  wire  [7:0] i_ifu_arlen,
    input  wire  [2:0] i_ifu_arsize,
    input  wire  [1:0] i_ifu_arburst,
    input  wire        i_ifu_arlock,
    input  wire  [3:0] i_ifu_arcache,
    input  wire  [2:0] i_ifu_arprot,
    input  wire  [3:0] i_ifu_arregion,
    input  wire  [3:0] i_ifu_arqos,
    input  wire        i_ifu_arvalid,
    output wire        o_ifu_arready,
    output wire  [2:0] o_ifu_rid,
    output wire [63:0] o_ifu_rdata,
    output wire  [1:0] o_ifu_rresp,
    output wire        o_ifu_rlast,
    output wire        o_ifu_rvalid,
    input  wire        i_ifu_rready,
    input  wire  [3:0] i_lsu_awid,
    input  wire [31:0] i_lsu_awaddr,
    input  wire  [7:0] i_lsu_awlen,
    input  wire  [2:0] i_lsu_awsize,
    input  wire  [1:0] i_lsu_awburst,
    input  wire        i_lsu_awlock,
    input  wire  [3:0] i_lsu_awcache,
    input  wire  [2:0] i_lsu_awprot,
    input  wire  [3:0] i_lsu_awregion,
    input  wire  [3:0] i_lsu_awqos,
    input  wire        i_lsu_awvalid,
    output wire        o_lsu_awready,
    input  wire  [3:0] i_lsu_arid,
    input  wire [31:0] i_lsu_araddr,
    input  wire  [7:0] i_lsu_arlen,
    input  wire  [2:0] i_lsu_arsize,
    input  wire  [1:0] i_lsu_arburst,
    input  wire        i_lsu_arlock,
    input  wire  [3:0] i_lsu_arcache,
    input  wire  [2:0] i_lsu_arprot,
    input  wire  [3:0] i_lsu_arregion,
    input  wire  [3:0] i_lsu_arqos,
    input  wire        i_lsu_arvalid,
    output wire        o_lsu_arready,
    input  wire [63:0] i_lsu_wdata,
    input  wire  [7:0] i_lsu_wstrb,
    input  wire        i_lsu_wlast,
    input  wire        i_lsu_wvalid,
    output wire        o_lsu_wready,
    output wire  [3:0] o_lsu_bid,
    output wire  [1:0] o_lsu_bresp,
    output wire        o_lsu_bvalid,
    input  wire        i_lsu_bready,
    output wire  [3:0] o_lsu_rid,
    output wire [63:0] o_lsu_rdata,
    output wire  [1:0] o_lsu_rresp,
    output wire        o_lsu_rlast,
    output wire        o_lsu_rvalid,
    input  wire        i_lsu_rready,
    input  wire  [0:0] i_sb_awid,
    input  wire [31:0] i_sb_awaddr,
    input  wire  [7:0] i_sb_awlen,
    input  wire  [2:0] i_sb_awsize,
    input  wire  [1:0] i_sb_awburst,
    input  wire        i_sb_awlock,
    input  wire  [3:0] i_sb_awcache,
    input  wire  [2:0] i_sb_awprot,
    input  wire  [3:0] i_sb_awregion,
    input  wire  [3:0] i_sb_awqos,
    input  wire        i_sb_awvalid,
    output wire        o_sb_awready,
    input  wire  [0:0] i_sb_arid,
    input  wire [31:0] i_sb_araddr,
    input  wire  [7:0] i_sb_arlen,
    input  wire  [2:0] i_sb_arsize,
    input  wire  [1:0] i_sb_arburst,
    input  wire        i_sb_arlock,
    input  wire  [3:0] i_sb_arcache,
    input  wire  [2:0] i_sb_arprot,
    input  wire  [3:0] i_sb_arregion,
    input  wire  [3:0] i_sb_arqos,
    input  wire        i_sb_arvalid,
    output wire        o_sb_arready,
    input  wire [63:0] i_sb_wdata,
    input  wire  [7:0] i_sb_wstrb,
    input  wire        i_sb_wlast,
    input  wire        i_sb_wvalid,
    output wire        o_sb_wready,
    output wire  [0:0] o_sb_bid,
    output wire  [1:0] o_sb_bresp,
    output wire        o_sb_bvalid,
    input  wire        i_sb_bready,
    output wire  [0:0] o_sb_rid,
    output wire [63:0] o_sb_rdata,
    output wire  [1:0] o_sb_rresp,
    output wire        o_sb_rlast,
    output wire        o_sb_rvalid,
    input  wire        i_sb_rready,
    output wire  [5:0] o_io_awid,
    output wire [31:0] o_io_awaddr,
    output wire  [7:0] o_io_awlen,
    output wire  [2:0] o_io_awsize,
    output wire  [1:0] o_io_awburst,
    output wire        o_io_awlock,
    output wire  [3:0] o_io_awcache,
    output wire  [2:0] o_io_awprot,
    output wire  [3:0] o_io_awregion,
    output wire  [3:0] o_io_awqos,
    output wire        o_io_awvalid,
    input  wire        i_io_awready,
    output wire  [5:0] o_io_arid,
    output wire [31:0] o_io_araddr,
    output wire  [7:0] o_io_arlen,
    output wire  [2:0] o_io_arsize,
    output wire  [1:0] o_io_arburst,
    output wire        o_io_arlock,
    output wire  [3:0] o_io_arcache,
    output wire  [2:0] o_io_arprot,
    output wire  [3:0] o_io_arregion,
    output wire  [3:0] o_io_arqos,
    output wire        o_io_arvalid,
    input  wire        i_io_arready,
    output wire [63:0] o_io_wdata,
    output wire  [7:0] o_io_wstrb,
    output wire        o_io_wlast,
    output wire        o_io_wvalid,
    input  wire        i_io_wready,
    input  wire  [5:0] i_io_bid,
    input  wire  [1:0] i_io_bresp,
    input  wire        i_io_bvalid,
    output wire        o_io_bready,
    input  wire  [5:0] i_io_rid,
    input  wire [63:0] i_io_rdata,
    input  wire  [1:0] i_io_rresp,
    input  wire        i_io_rlast,
    input  wire        i_io_rvalid,
    output wire        o_io_rready,
    output wire  [5:0] o_ram_awid,
    output wire [31:0] o_ram_awaddr,
    output wire  [7:0] o_ram_awlen,
    output wire  [2:0] o_ram_awsize,
    output wire  [1:0] o_ram_awburst,
    output wire        o_ram_awlock,
    output wire  [3:0] o_ram_awcache,
    output wire  [2:0] o_ram_awprot,
    output wire  [3:0] o_ram_awregion,
    output wire  [3:0] o_ram_awqos,
    output wire        o_ram_awvalid,
    input  wire        i_ram_awready,
    output wire  [5:0] o_ram_arid,
    output wire [31:0] o_ram_araddr,
    output wire  [7:0] o_ram_arlen,
    output wire  [2:0] o_ram_arsize,
    output wire  [1:0] o_ram_arburst,
    output wire        o_ram_arlock,
    output wire  [3:0] o_ram_arcache,
    output wire  [2:0] o_ram_arprot,
    output wire  [3:0] o_ram_arregion,
    output wire  [3:0] o_ram_arqos,
    output wire        o_ram_arvalid,
    input  wire        i_ram_arready,
    output wire [63:0] o_ram_wdata,
    output wire  [7:0] o_ram_wstrb,
    output wire        o_ram_wlast,
    output wire        o_ram_wvalid,
    input  wire        i_ram_wready,
    input  wire  [5:0] i_ram_bid,
    input  wire  [1:0] i_ram_bresp,
    input  wire        i_ram_bvalid,
    output wire        o_ram_bready,
    input  wire  [5:0] i_ram_rid,
    input  wire [63:0] i_ram_rdata,
    input  wire  [1:0] i_ram_rresp,
    input  wire        i_ram_rlast,
    input  wire        i_ram_rvalid,
    output wire        o_ram_rready,
	
	output wire  [5:0] o_user_awid,
    output wire [31:0] o_user_awaddr,
    output wire  [7:0] o_user_awlen,
    output wire  [2:0] o_user_awsize,
    output wire  [1:0] o_user_awburst,
    output wire        o_user_awlock,
    output wire  [3:0] o_user_awcache,
    output wire  [2:0] o_user_awprot,
    output wire  [3:0] o_user_awregion,
    output wire  [3:0] o_user_awqos,
    output wire        o_user_awvalid,
    input  wire        i_user_awready,
    output wire  [5:0] o_user_arid,
    output wire [31:0] o_user_araddr,
    output wire  [7:0] o_user_arlen,
    output wire  [2:0] o_user_arsize,
    output wire  [1:0] o_user_arburst,
    output wire        o_user_arlock,
    output wire  [3:0] o_user_arcache,
    output wire  [2:0] o_user_arprot,
    output wire  [3:0] o_user_arregion,
    output wire  [3:0] o_user_arqos,
    output wire        o_user_arvalid,
    input  wire        i_user_arready,
    output wire [63:0] o_user_wdata,
    output wire  [7:0] o_user_wstrb,
    output wire        o_user_wlast,
    output wire        o_user_wvalid,
    input  wire        i_user_wready,
    input  wire  [5:0] i_user_bid,
    input  wire  [1:0] i_user_bresp,
    input  wire        i_user_bvalid,
    output wire        o_user_bready,
    input  wire  [5:0] i_user_rid,
    input  wire [63:0] i_user_rdata,
    input  wire  [1:0] i_user_rresp,
    input  wire        i_user_rlast,
    input  wire        i_user_rvalid,
    output wire        o_user_rready
);
 
axi_intercon axi_intercon2
   (
    .clk_i              (clk_i),
    .rst_ni             (rst_ni),
    .i_ifu_arid         (i_ifu_arid),
    .i_ifu_araddr       (i_ifu_araddr),
    .i_ifu_arlen        (i_ifu_arlen),
    .i_ifu_arsize       (i_ifu_arsize),
    .i_ifu_arburst      (i_ifu_arburst),
    .i_ifu_arlock       (i_ifu_arlock),
    .i_ifu_arcache      (i_ifu_arcache),
    .i_ifu_arprot       (i_ifu_arprot),
    .i_ifu_arregion     (i_ifu_arregion),
    .i_ifu_arqos        (i_ifu_arqos),
    .i_ifu_arvalid      (i_ifu_arvalid),
    .o_ifu_arready      (o_ifu_arready),
    .o_ifu_rid          (o_ifu_rid),
    .o_ifu_rdata        (o_ifu_rdata),
    .o_ifu_rresp        (o_ifu_rresp),
    .o_ifu_rlast        (o_ifu_rlast),
    .o_ifu_rvalid       (o_ifu_rvalid),
    .i_ifu_rready       (i_ifu_rready),
    .i_lsu_awid         (i_lsu_awid),
    .i_lsu_awaddr       (i_lsu_awaddr),
    .i_lsu_awlen        (i_lsu_awlen),
    .i_lsu_awsize       (i_lsu_awsize),
    .i_lsu_awburst      (i_lsu_awburst),
    .i_lsu_awlock       (i_lsu_awlock),  
    .i_lsu_awcache      (i_lsu_awcache),
    .i_lsu_awprot       (i_lsu_awprot),
    .i_lsu_awregion     (i_lsu_awregion),
    .i_lsu_awqos        (i_lsu_awqos),
    .i_lsu_awvalid      (i_lsu_awvalid),
    .o_lsu_awready      (o_lsu_awready),
    .i_lsu_arid         (i_lsu_arid),
    .i_lsu_araddr       (i_lsu_araddr),
    .i_lsu_arlen        (i_lsu_arlen),
    .i_lsu_arsize       (i_lsu_arsize),
    .i_lsu_arburst      (i_lsu_arburst),
    .i_lsu_arlock       (i_lsu_arlock),
    .i_lsu_arcache      (i_lsu_arcache),
    .i_lsu_arprot       (i_lsu_arprot),
    .i_lsu_arregion     (i_lsu_arregion),
    .i_lsu_arqos        (i_lsu_arqos),
    .i_lsu_arvalid      (i_lsu_arvalid),
    .o_lsu_arready      (o_lsu_arready),
    .i_lsu_wdata        (i_lsu_wdata),
    .i_lsu_wstrb        (i_lsu_wstrb),
    .i_lsu_wlast        (i_lsu_wlast),
    .i_lsu_wvalid       (i_lsu_wvalid),
    .o_lsu_wready       (o_lsu_wready),
    .o_lsu_bid          (o_lsu_bid),
    .o_lsu_bresp        (o_lsu_bresp),
    .o_lsu_bvalid       (o_lsu_bvalid),
    .i_lsu_bready       (i_lsu_bready),
    .o_lsu_rid          (o_lsu_rid),
    .o_lsu_rdata        (o_lsu_rdata),
    .o_lsu_rresp        (o_lsu_rresp),
    .o_lsu_rlast        (o_lsu_rlast),
    .o_lsu_rvalid       (o_lsu_rvalid),
    .i_lsu_rready       (i_lsu_rready),
    .i_sb_awid          (i_sb_awid),
    .i_sb_awaddr        (i_sb_awaddr),
    .i_sb_awlen         (i_sb_awlen),
    .i_sb_awsize        (i_sb_awsize),
    .i_sb_awburst       (i_sb_awburst),
    .i_sb_awlock        (i_sb_awlock),
    .i_sb_awcache       (i_sb_awcache),
    .i_sb_awprot        (i_sb_awprot),
    .i_sb_awregion      (i_sb_awregion),
    .i_sb_awqos         (i_sb_awqos),
    .i_sb_awvalid       (i_sb_awvalid),
    .o_sb_awready       (o_sb_awready),
    .i_sb_arid          (i_sb_arid),
    .i_sb_araddr        (i_sb_araddr),
    .i_sb_arlen         (i_sb_arlen),
    .i_sb_arsize        (i_sb_arsize),
    .i_sb_arburst       (i_sb_arburst),
    .i_sb_arlock        (i_sb_arlock),
    .i_sb_arcache       (i_sb_arcache),
    .i_sb_arprot        (i_sb_arprot),
    .i_sb_arregion      (i_sb_arregion),
    .i_sb_arqos         (i_sb_arqos),
    .i_sb_arvalid       (i_sb_arvalid),
    .o_sb_arready       (o_sb_arready),
    .i_sb_wdata         (i_sb_wdata),
    .i_sb_wstrb         (i_sb_wstrb),
    .i_sb_wlast         (i_sb_wlast),
    .i_sb_wvalid        (i_sb_wvalid),
    .o_sb_wready        (o_sb_wready),
    .o_sb_bid           (o_sb_bid),
    .o_sb_bresp         (o_sb_bresp),
    .o_sb_bvalid        (o_sb_bvalid),
    .i_sb_bready        (i_sb_bready),
    .o_sb_rid           (o_sb_rid),
    .o_sb_rdata         (o_sb_rdata),
    .o_sb_rresp         (o_sb_rresp),
    .o_sb_rlast         (o_sb_rlast),
    .o_sb_rvalid        (o_sb_rvalid),
    .i_sb_rready        (i_sb_rready),
    .o_io_awid          (o_io_awid),
    .o_io_awaddr        (o_io_awaddr),
    .o_io_awlen         (o_io_awlen),
    .o_io_awsize        (o_io_awsize),
    .o_io_awburst       (o_io_awburst),
    .o_io_awlock        (o_io_awlock),
    .o_io_awcache       (o_io_awcache),
    .o_io_awprot        (o_io_awprot),
    .o_io_awregion      (o_io_awregion),
    .o_io_awqos         (o_io_awqos),
    .o_io_awvalid       (o_io_awvalid),
    .i_io_awready       (i_io_awready),
    .o_io_arid          (o_io_arid),
    .o_io_araddr        (o_io_araddr),
    .o_io_arlen         (o_io_arlen),
    .o_io_arsize        (o_io_arsize),
    .o_io_arburst       (o_io_arburst),
    .o_io_arlock        (o_io_arlock),
    .o_io_arcache       (o_io_arcache),
    .o_io_arprot        (o_io_arprot),
    .o_io_arregion      (o_io_arregion),
    .o_io_arqos         (o_io_arqos),
    .o_io_arvalid       (o_io_arvalid),
    .i_io_arready       (i_io_arready),
    .o_io_wdata         (o_io_wdata),
    .o_io_wstrb         (o_io_wstrb),
    .o_io_wlast         (o_io_wlast),
    .o_io_wvalid        (o_io_wvalid),
    .i_io_wready        (i_io_wready),
    .i_io_bid           (i_io_bid),
    .i_io_bresp         (i_io_bresp),
    .i_io_bvalid        (i_io_bvalid),
    .o_io_bready        (o_io_bready),
    .i_io_rid           (i_io_rid),
    .i_io_rdata         (i_io_rdata),
    .i_io_rresp         (i_io_rresp),
    .i_io_rlast         (i_io_rlast),
    .i_io_rvalid        (i_io_rvalid),
    .o_io_rready        (o_io_rready),
    .o_ram_awid         (o_ram_awid),
    .o_ram_awaddr       (o_ram_awaddr),
    .o_ram_awlen        (o_ram_awlen),
    .o_ram_awsize       (o_ram_awsize),
    .o_ram_awburst       (o_ram_awburst),
    .o_ram_awlock       (o_ram_awlock),
    .o_ram_awcache      (o_ram_awcache),
    .o_ram_awprot       (o_ram_awprot),
    .o_ram_awregion     (o_ram_awregion),
    .o_ram_awqos        (o_ram_awqos),
    .o_ram_awvalid      (o_ram_awvalid),
    .i_ram_awready      (i_ram_awready),
    .o_ram_arid         (o_ram_arid),
    .o_ram_araddr       (o_ram_araddr),
    .o_ram_arlen        (o_ram_arlen),
    .o_ram_arsize       (o_ram_arsize),
    .o_ram_arburst      (o_ram_arburst),
    .o_ram_arlock       (o_ram_arlock),
    .o_ram_arcache      (o_ram_arcache),
    .o_ram_arprot       (o_ram_arprot),
    .o_ram_arregion     (o_ram_arregion),
    .o_ram_arqos        (o_ram_arqos),
    .o_ram_arvalid      (o_ram_arvalid),
    .i_ram_arready      (i_ram_arready),
    .o_ram_wdata        (o_ram_wdata),
    .o_ram_wstrb        (o_ram_wstrb),
    .o_ram_wlast        (o_ram_wlast),
    .o_ram_wvalid       (o_ram_wvalid),
    .i_ram_wready       (i_ram_wready),
    .i_ram_bid          (i_ram_bid),
    .i_ram_bresp        (i_ram_bresp),
    .i_ram_bvalid       (i_ram_bvalid),
    .o_ram_bready       (o_ram_bready),
    .i_ram_rid          (i_ram_rid),
    .i_ram_rdata        (i_ram_rdata),
    .i_ram_rresp        (i_ram_rresp),
    .i_ram_rlast        (i_ram_rlast),
    .i_ram_rvalid       (i_ram_rvalid),
    .o_ram_rready       (o_ram_rready),
	.o_user_awid		(o_user_awid),
	.o_user_awaddr		(o_user_awaddr),
	.o_user_awlen		(o_user_awlen),
	.o_user_awsize		(o_user_awsize),
	.o_user_awburst		(o_user_awburst),
	.o_user_awlock		(o_user_awlock),
	.o_user_awcache		(o_user_awcache),
	.o_user_awprot		(o_user_awprot),
	.o_user_awregion	(o_user_awregion),
	.o_user_awqos		(o_user_awqos),
	.o_user_awvalid		(o_user_awvalid),
	.i_user_awready		(i_user_awready),
	.o_user_arid		(o_user_arid),
	.o_user_araddr		(o_user_araddr),
	.o_user_arlen		(o_user_arlen),
	.o_user_arsize		(o_user_arsize),
	.o_user_arburst		(o_user_arburst),
	.o_user_arlock		(o_user_arlock),
	.o_user_arcache		(o_user_arcache),
	.o_user_arprot		(o_user_arprot),
	.o_user_arregion	(o_user_arregion),
	.o_user_arqos		(o_user_arqos),
	.o_user_arvalid		(o_user_arvalid),
	.i_user_arready		(i_user_arready),
	.o_user_wdata		(o_user_wdata),
	.o_user_wstrb		(o_user_wstrb),
	.o_user_wlast		(o_user_wlast),
	.o_user_wvalid		(o_user_wvalid),
	.i_user_wready		(i_user_wready),
	.i_user_bid			(i_user_bid),
	.i_user_bresp		(i_user_bresp),
	.i_user_bvalid		(i_user_bvalid),
	.o_user_bready		(o_user_bready),
	.i_user_rid			(i_user_rid),
	.i_user_rdata		(i_user_rdata),
	.i_user_rresp		(i_user_rresp),
	.i_user_rlast		(i_user_rlast),
	.i_user_rvalid		(i_user_rvalid),
	.o_user_rready		(o_user_rready)
    );
    
endmodule


